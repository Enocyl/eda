`timescale 1ns / 1ns
// `default_nettype none

// 80bit output 0

module const_0_80b (dout);

    output [79:0] dout;


    // dout  80bit
    assign dout = 80'd0;

endmodule