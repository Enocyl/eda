module buf8b(I, 
             O);

    input [7:0] I;
   output [7:0] O;
   
   
   BUF  XLXI_1 (.I(I[0]), 
               .O(O[0]));
   BUF  XLXI_2 (.I(I[1]), 
               .O(O[1]));
   BUF  XLXI_3 (.I(I[2]), 
               .O(O[2]));
   BUF  XLXI_4 (.I(I[3]), 
               .O(O[3]));
   BUF  XLXI_5 (.I(I[4]), 
               .O(O[4]));
   BUF  XLXI_6 (.I(I[5]), 
               .O(O[5]));
   BUF  XLXI_7 (.I(I[6]), 
               .O(O[6]));
   BUF  XLXI_8 (.I(I[7]), 
               .O(O[7]));
endmodule
