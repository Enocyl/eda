module m8_1e16b(E, 
                                    I0D, 
                                    I1D, 
                                    I2D, 
                                    I3D, 
                                    I4D, 
                                    I5D, 
                                    I6D, 
                                    I7D, 
                                    S, 
                                    O);

    input E;
    input [15:0] I0D;
    input [15:0] I1D;
    input [15:0] I2D;
    input [15:0] I3D;
    input [15:0] I4D;
    input [15:0] I5D;
    input [15:0] I6D;
    input [15:0] I7D;
    input [2:0] S;
   output [15:0] O;
   
   
   (* HU_SET = "XLXI_73_9" *) 
   M8_1E  XLXI_73 (.D0(I0D[0]), 
                                        .D1(I1D[0]), 
                                        .D2(I2D[0]), 
                                        .D3(I3D[0]), 
                                        .D4(I4D[0]), 
                                        .D5(I5D[0]), 
                                        .D6(I6D[0]), 
                                        .D7(I7D[0]), 
                                        .E(E), 
                                        .S0(S[0]), 
                                        .S1(S[1]), 
                                        .S2(S[2]), 
                                        .O(O[0]));
   (* HU_SET = "XLXI_74_10" *) 
   M8_1E  XLXI_74 (.D0(I0D[1]), 
                                        .D1(I1D[1]), 
                                        .D2(I2D[1]), 
                                        .D3(I3D[1]), 
                                        .D4(I4D[1]), 
                                        .D5(I5D[1]), 
                                        .D6(I6D[1]), 
                                        .D7(I7D[1]), 
                                        .E(E), 
                                        .S0(S[0]), 
                                        .S1(S[1]), 
                                        .S2(S[2]), 
                                        .O(O[1]));
   (* HU_SET = "XLXI_75_12" *) 
   M8_1E  XLXI_75 (.D0(I0D[3]), 
                                        .D1(I1D[3]), 
                                        .D2(I2D[3]), 
                                        .D3(I3D[3]), 
                                        .D4(I4D[3]), 
                                        .D5(I5D[3]), 
                                        .D6(I6D[3]), 
                                        .D7(I7D[3]), 
                                        .E(E), 
                                        .S0(S[0]), 
                                        .S1(S[1]), 
                                        .S2(S[2]), 
                                        .O(O[3]));
   (* HU_SET = "XLXI_76_11" *) 
   M8_1E  XLXI_76 (.D0(I0D[2]), 
                                        .D1(I1D[2]), 
                                        .D2(I2D[2]), 
                                        .D3(I3D[2]), 
                                        .D4(I4D[2]), 
                                        .D5(I5D[2]), 
                                        .D6(I6D[2]), 
                                        .D7(I7D[2]), 
                                        .E(E), 
                                        .S0(S[0]), 
                                        .S1(S[1]), 
                                        .S2(S[2]), 
                                        .O(O[2]));
   (* HU_SET = "XLXI_77_13" *) 
   M8_1E  XLXI_77 (.D0(I0D[4]), 
                                        .D1(I1D[4]), 
                                        .D2(I2D[4]), 
                                        .D3(I3D[4]), 
                                        .D4(I4D[4]), 
                                        .D5(I5D[4]), 
                                        .D6(I6D[4]), 
                                        .D7(I7D[4]), 
                                        .E(E), 
                                        .S0(S[0]), 
                                        .S1(S[1]), 
                                        .S2(S[2]), 
                                        .O(O[4]));
   (* HU_SET = "XLXI_78_14" *) 
   M8_1E  XLXI_78 (.D0(I0D[5]), 
                                        .D1(I1D[5]), 
                                        .D2(I2D[5]), 
                                        .D3(I3D[5]), 
                                        .D4(I4D[5]), 
                                        .D5(I5D[5]), 
                                        .D6(I6D[5]), 
                                        .D7(I7D[5]), 
                                        .E(E), 
                                        .S0(S[0]), 
                                        .S1(S[1]), 
                                        .S2(S[2]), 
                                        .O(O[5]));
   (* HU_SET = "XLXI_79_16" *) 
   M8_1E  XLXI_79 (.D0(I0D[7]), 
                                        .D1(I1D[7]), 
                                        .D2(I2D[7]), 
                                        .D3(I3D[7]), 
                                        .D4(I4D[7]), 
                                        .D5(I5D[7]), 
                                        .D6(I6D[7]), 
                                        .D7(I7D[7]), 
                                        .E(E), 
                                        .S0(S[0]), 
                                        .S1(S[1]), 
                                        .S2(S[2]), 
                                        .O(O[7]));
   (* HU_SET = "XLXI_80_15" *) 
   M8_1E  XLXI_80 (.D0(I0D[6]), 
                                        .D1(I1D[6]), 
                                        .D2(I2D[6]), 
                                        .D3(I3D[6]), 
                                        .D4(I4D[6]), 
                                        .D5(I5D[6]), 
                                        .D6(I6D[6]), 
                                        .D7(I7D[6]), 
                                        .E(E), 
                                        .S0(S[0]), 
                                        .S1(S[1]), 
                                        .S2(S[2]), 
                                        .O(O[6]));
   (* HU_SET = "XLXI_81_17" *) 
   M8_1E  XLXI_81 (.D0(I0D[8]), 
                                        .D1(I1D[8]), 
                                        .D2(I2D[8]), 
                                        .D3(I3D[8]), 
                                        .D4(I4D[8]), 
                                        .D5(I5D[8]), 
                                        .D6(I6D[8]), 
                                        .D7(I7D[8]), 
                                        .E(E), 
                                        .S0(S[0]), 
                                        .S1(S[1]), 
                                        .S2(S[2]), 
                                        .O(O[8]));
   (* HU_SET = "XLXI_82_18" *) 
   M8_1E  XLXI_82 (.D0(I0D[9]), 
                                        .D1(I1D[9]), 
                                        .D2(I2D[9]), 
                                        .D3(I3D[9]), 
                                        .D4(I4D[9]), 
                                        .D5(I5D[9]), 
                                        .D6(I6D[9]), 
                                        .D7(I7D[9]), 
                                        .E(E), 
                                        .S0(S[0]), 
                                        .S1(S[1]), 
                                        .S2(S[2]), 
                                        .O(O[9]));
   (* HU_SET = "XLXI_118_19" *) 
   M8_1E  XLXI_118 (.D0(I0D[10]), 
                                         .D1(I1D[10]), 
                                         .D2(I2D[10]), 
                                         .D3(I3D[10]), 
                                         .D4(I4D[10]), 
                                         .D5(I5D[10]), 
                                         .D6(I6D[10]), 
                                         .D7(I7D[10]), 
                                         .E(E), 
                                         .S0(S[0]), 
                                         .S1(S[1]), 
                                         .S2(S[2]), 
                                         .O(O[10]));
   (* HU_SET = "XLXI_119_20" *) 
   M8_1E  XLXI_119 (.D0(I0D[11]), 
                                         .D1(I1D[11]), 
                                         .D2(I2D[11]), 
                                         .D3(I3D[11]), 
                                         .D4(I4D[11]), 
                                         .D5(I5D[11]), 
                                         .D6(I6D[11]), 
                                         .D7(I7D[11]), 
                                         .E(E), 
                                         .S0(S[0]), 
                                         .S1(S[1]), 
                                         .S2(S[2]), 
                                         .O(O[11]));
   (* HU_SET = "XLXI_144_21" *) 
   M8_1E  XLXI_144 (.D0(I0D[12]), 
                                         .D1(I1D[12]), 
                                         .D2(I2D[12]), 
                                         .D3(I3D[12]), 
                                         .D4(I4D[12]), 
                                         .D5(I5D[12]), 
                                         .D6(I6D[12]), 
                                         .D7(I7D[12]), 
                                         .E(E), 
                                         .S0(S[0]), 
                                         .S1(S[1]), 
                                         .S2(S[2]), 
                                         .O(O[12]));
   (* HU_SET = "XLXI_145_22" *) 
   M8_1E  XLXI_145 (.D0(I0D[13]), 
                                         .D1(I1D[13]), 
                                         .D2(I2D[13]), 
                                         .D3(I3D[13]), 
                                         .D4(I4D[13]), 
                                         .D5(I5D[13]), 
                                         .D6(I6D[13]), 
                                         .D7(I7D[13]), 
                                         .E(E), 
                                         .S0(S[0]), 
                                         .S1(S[1]), 
                                         .S2(S[2]), 
                                         .O(O[13]));
   (* HU_SET = "XLXI_146_23" *) 
   M8_1E  XLXI_146 (.D0(I0D[14]), 
                                         .D1(I1D[14]), 
                                         .D2(I2D[14]), 
                                         .D3(I3D[14]), 
                                         .D4(I4D[14]), 
                                         .D5(I5D[14]), 
                                         .D6(I6D[14]), 
                                         .D7(I7D[14]), 
                                         .E(E), 
                                         .S0(S[0]), 
                                         .S1(S[1]), 
                                         .S2(S[2]), 
                                         .O(O[14]));
   (* HU_SET = "XLXI_147_24" *) 
   M8_1E  XLXI_147 (.D0(I0D[15]), 
                                         .D1(I1D[15]), 
                                         .D2(I2D[15]), 
                                         .D3(I3D[15]), 
                                         .D4(I4D[15]), 
                                         .D5(I5D[15]), 
                                         .D6(I6D[15]), 
                                         .D7(I7D[15]), 
                                         .E(E), 
                                         .S0(S[0]), 
                                         .S1(S[1]), 
                                         .S2(S[2]), 
                                         .O(O[15]));
endmodule